package axi_enum;
// might needed enums
// enum for AXI states
// AXI states for read and write channels
//axi handshake states

endpackage 