package axi_constraints;
// Class:AXI constraints read package
//Class:AXI Constraints write package
//Class:AXI constraints for handshake signals
//Class:AXI constraints for memory 
endpackage